// Copyright 2020 ETH Zurich and University of Bologna.
// All rights reserved.
//
// This code is under development and not yet released to the public.
// Until it is released, the code is under the copyright of ETH Zurich and
// the University of Bologna, and may contain confidential and/or unpublished
// work. Any reuse/redistribution is strictly forbidden without written
// permission from ETH Zurich.

package automatic pspin_tb_cfg_pkg;
  // TB Parameters
  parameter time          CLK_PERIOD = 1000ps;

  //Debug
  parameter int unsigned  Verbosity = 0;

endpackage